/**
 *  bsg_cache_miss.v
 *
 *  miss handling unit.
 *
 *  @author tommy
 *
 */

`include "bsg_defines.v"
`include "bsg_cache.vh"

module bsg_cache_miss
  import bsg_cache_pkg::*;
  #(parameter `BSG_INV_PARAM(addr_width_p)
    ,parameter `BSG_INV_PARAM(data_width_p)
    ,parameter `BSG_INV_PARAM(block_size_in_words_p)
    ,parameter `BSG_INV_PARAM(sets_p)
    ,parameter `BSG_INV_PARAM(ways_p)
    ,parameter `BSG_INV_PARAM(word_tracking_p)

    ,parameter lg_block_size_in_words_lp=`BSG_SAFE_CLOG2(block_size_in_words_p)
    ,parameter lg_sets_lp=`BSG_SAFE_CLOG2(sets_p)
    ,parameter data_mask_width_lp=(data_width_p>>3)
    ,parameter lg_data_mask_width_lp=`BSG_SAFE_CLOG2(data_width_p>>3)
    ,parameter block_offset_width_lp=(block_size_in_words_p > 1) ? lg_data_mask_width_lp+lg_block_size_in_words_lp : lg_data_mask_width_lp
    ,parameter tag_width_lp=(addr_width_p-lg_sets_lp-block_offset_width_lp)
    ,parameter tag_info_width_lp=`bsg_cache_tag_info_width(tag_width_lp)
    ,parameter lg_ways_lp=`BSG_SAFE_CLOG2(ways_p)
    ,parameter stat_info_width_lp=`bsg_cache_stat_info_width(ways_p)
  )
  (
    input clk_i
    ,input reset_i

    // from tv stage
    ,input miss_v_i
    ,input track_miss_i
    ,input bsg_cache_decode_s decode_v_i
    ,input [addr_width_p-1:0] addr_v_i
    ,input [data_mask_width_lp-1:0] mask_v_i
    
    ,input [ways_p-1:0][tag_width_lp-1:0] tag_v_i
    ,input [ways_p-1:0] valid_v_i
    ,input [ways_p-1:0] lock_v_i
    ,input [ways_p-1:0] tag_hit_v_i

    ,input [lg_ways_lp-1:0] tag_hit_way_id_i
    ,input tag_hit_found_i
    ,input [data_width_p-1:0] data_v_i 

    // from store buffer
    ,input sbuf_empty_i

    // from track buffer
    ,input tbuf_empty_i

    // to dma engine
    ,output bsg_cache_dma_cmd_e         dma_cmd_o
    ,output logic [lg_ways_lp-1:0]      dma_way_o
    ,output logic [addr_width_p-1:0]    dma_addr_o
    ,input                              dma_done_i

    // to dma engine for flopping track_mem's read data
    // used to avoid clk-to-q timing from memory
    ,output logic track_data_we_o

    // from stat_mem
    ,input [stat_info_width_lp-1:0] stat_info_i

    // to stat_mem
    ,output logic stat_mem_v_o
    ,output logic stat_mem_w_o
    ,output logic [lg_sets_lp-1:0] stat_mem_addr_o
    ,output logic [stat_info_width_lp-1:0] stat_mem_data_o
    ,output logic [stat_info_width_lp-1:0] stat_mem_w_mask_o

    // to tag_mem
    ,output logic tag_mem_v_o
    ,output logic tag_mem_w_o
    ,output logic [lg_sets_lp-1:0] tag_mem_addr_o
    ,output logic [ways_p-1:0][tag_info_width_lp-1:0] tag_mem_data_o
    ,output logic [ways_p-1:0][tag_info_width_lp-1:0] tag_mem_w_mask_o

    // to track mem
    ,output logic track_mem_v_o
    ,output logic track_mem_w_o
    ,output logic [lg_sets_lp-1:0] track_mem_addr_o
    ,output logic [ways_p-1:0][block_size_in_words_p-1:0] track_mem_w_mask_o
    ,output logic [ways_p-1:0][block_size_in_words_p-1:0] track_mem_data_o

    // to pipeline
    ,output logic                                 done_o
    ,output logic                                 recover_o
    ,output logic [lg_ways_lp-1:0]                chosen_way_o
    ,output logic                                 select_snoop_data_r_o
    ,output logic                                 miss_active_o
    ,output logic                                 dma_stall_o
    ,output logic                                 id
    ,output [data_width_p-1:0]                    data_o

    ,output logic [data_mask_width_lp-1:0]        mask_v_miss_o
    ,output bsg_cache_decode_s                    decode_v_miss_o
    ,output logic [tag_width_lp-1:0]              addr_v_miss_o
    ,output logic [data_width_p-1:0]              data_v_miss_o
    ,output logic [ways_p-1:0]                    valid_v_miss_o
    ,output logic [ways_p-1:0][tag_width_lp-1:0]  tag_v_miss_o
    ,output logic [ways_p-1:0]                    lock_v_miss_o

    ,input ack_i
  );

  // stat/tag info
  //
  `declare_bsg_cache_tag_info_s(tag_width_lp);
  `declare_bsg_cache_stat_info_s(ways_p);

  bsg_cache_stat_info_s stat_info_in;
  assign stat_info_in = stat_info_i;

  bsg_cache_tag_info_s [ways_p-1:0] tag_mem_data_out, tag_mem_w_mask_out;
  bsg_cache_stat_info_s stat_mem_data_out, stat_mem_w_mask_out;
  
  assign tag_mem_data_o = tag_mem_data_out;
  assign stat_mem_data_o = stat_mem_data_out;

  assign tag_mem_w_mask_o = tag_mem_w_mask_out;
  assign stat_mem_w_mask_o = stat_mem_w_mask_out;


  // miss handler FSM
  //
  typedef enum logic [3:0] {
    START
    ,FLUSH_OP
    ,LOCK_OP
    ,SEND_EVICT_ADDR
    ,SEND_FILL_ADDR
    ,SEND_EVICT_DATA
    ,GET_FILL_DATA
    ,WAIT_FOR_FILL_DATA
    ,STORE_TAG_MISS
    ,STORE_TAG_MISS_ALLOCATE
    ,RECOVER
    ,DONE
  } miss_state_e;

  miss_state_e miss_state_r;
  miss_state_e miss_state_n;
  logic [lg_ways_lp-1:0] chosen_way_r, chosen_way_n;
  logic [lg_ways_lp-1:0] flush_way_r, flush_way_n;
  logic select_snoop_data_r, select_snoop_data_n;

  logic [tag_width_lp-1:0] addr_tag_v;
  logic [lg_sets_lp-1:0] addr_index_v;
  logic [lg_ways_lp-1:0] addr_way_v;
  logic [lg_block_size_in_words_lp-1:0] addr_block_offset_v;

  // for flush/inv ops, go to FLUSH_OP.
  // for AUNLOCK, or ALOCK with tag hit, to go LOCK_OP.
  // for store tag miss with data size equal or bigger than a word, do not fetch cache line word tracking is enables

  wire goto_flush_op = decode_v_i.tagfl_op| decode_v_i.ainv_op| decode_v_i.afl_op| decode_v_i.aflinv_op;
  wire goto_lock_op = decode_v_i.aunlock_op | (decode_v_i.alock_op & tag_hit_found_i);
  wire full_word_op = decode_v_i.mask_op
    ? (&mask_v_i)
    : (decode_v_i.data_size_op >= lg_data_mask_width_lp);
  wire st_tag_miss_op = word_tracking_p ? (decode_v_i.st_op & full_word_op & ~tag_hit_found_i) : 1'b0;
 
  logic [data_mask_width_lp-1:0]        mask_v_r;
  bsg_cache_decode_s                    decode_v_r;
  logic [tag_width_lp-1:0]              addr_tag_v_r;
  logic [lg_sets_lp-1:0]                addr_index_v_r;
  logic [lg_ways_lp-1:0]                addr_way_v_r;
  logic [lg_block_size_in_words_lp-1:0] addr_block_offset_v_r;
  logic [data_width_p-1:0]              data_v_r;
  logic [ways_p-1:0]                    valid_v_r;
  logic [ways_p-1:0][tag_width_lp-1:0]  tag_v_r;
  logic [ways_p-1:0]                    lock_v_r;

  logic [ways_p-1:0]                    tag_hit_v_r;
  logic [lg_ways_lp-1:0]                tag_hit_way_id_r;
  logic                                 tag_hit_found_r;

  logic goto_flush_op_r;
  logic goto_lock_op_r;
  logic st_tag_miss_op_r;
  logic track_miss_r;
  logic [addr_width_p-1:0] addr_v_r;
   
  // Capture all information from tag verify stage for miss handling
  // Capture when there is a valid miss and not when the state machine is
  // active
  always_ff @(posedge clk_i) begin
    if(miss_v_i & ~miss_active_o) begin
      addr_v_r              <= addr_v_i;
      data_v_r              <= data_v_i;
      track_miss_r          <= track_miss_i;
      tag_v_r               <= tag_v_i;
      tag_hit_v_r           <= tag_hit_v_i;
      lock_v_r              <= lock_v_i;
      tag_hit_way_id_r      <= tag_hit_way_id_i;
      tag_hit_found_r       <= tag_hit_found_i;
      decode_v_r            <= decode_v_i;
      mask_v_r              <= mask_v_i;
      valid_v_r             <= valid_v_i;
      goto_flush_op_r       <= goto_flush_op;
      goto_lock_op_r        <= goto_lock_op;
      st_tag_miss_op_r      <= st_tag_miss_op;
    end
  end
  
  assign addr_index_v_r           = addr_v_r[block_offset_width_lp+:lg_sets_lp];
  assign addr_tag_v_r             = addr_v_r[block_offset_width_lp+lg_sets_lp+:tag_width_lp];
  assign addr_way_v_r             = addr_v_r[block_offset_width_lp+lg_sets_lp+:lg_ways_lp];
  assign addr_block_offset_v_r    = addr_v_r[lg_data_mask_width_lp+:lg_block_size_in_words_lp];

  assign mask_v_miss_o          = mask_v_r;
  assign decode_v_miss_o        = decode_v_r;
  assign addr_v_miss_o          = addr_v_r;
  assign data_v_miss_o          = data_v_r;
  assign valid_v_miss_o         = valid_v_r;
  assign tag_v_miss_o           = tag_v_r;
  assign lock_v_miss_o          = lock_v_r;

    
  // Check if address match from tl stage and send data
  //always_comb begin 
  //  tag_tl_hit = 1'b0;
  //  if((addr_tag_tl == addr_tag_v_r) && (addr_index_tl == addr_index_v_r)) begin 
  //      tag_tl_hit = 1'b1;
  //  end
  //end
  
  // Communicate to the pipeline that a miss is currently being serviced
  assign miss_active_o = (miss_state_r != START);
  assign id = miss_active_o & (miss_state_r != DONE);
  
  // Find the way that is invalid.
  //
  logic [lg_ways_lp-1:0] invalid_way_id;
  logic invalid_exist;

  bsg_priority_encode #(
    .width_p(ways_p)
    ,.lo_to_hi_p(1)
  ) invalid_way_pe (
    .i(~valid_v_r & ~lock_v_r) // invalid and unlocked
    ,.addr_o(invalid_way_id)
    ,.v_o(invalid_exist)
  );

  assign stat_mem_addr_o = addr_index_v_r;
  assign tag_mem_addr_o = addr_index_v_r;
  assign track_mem_addr_o = addr_index_v_r;

  assign chosen_way_o = chosen_way_r;

  assign dma_way_o = goto_flush_op_r
    ? flush_way_r
    : chosen_way_r;

  // chosen way lru decode
  //
  logic [ways_p-2:0] chosen_way_lru_data;
  logic [ways_p-2:0] chosen_way_lru_mask;

  bsg_lru_pseudo_tree_decode #(
    .ways_p(ways_p)
  ) chosen_way_lru_decode (
    .way_id_i(chosen_way_r)
    ,.data_o(chosen_way_lru_data)
    ,.mask_o(chosen_way_lru_mask)
  );

  // backup LRU
  // When the LRU way designated by the stats_mem_info is locked, a backup way is required for 
  // cache line replacement. In the current design, bsg_lru_pseudo_tree_backup takes the way with 
  // the shortest distance from the locked LRU way in the tree, as the backup option by overriding
  // some of the LRU bits, so that it avoids "LRU trap" from insufficient update on the LRU bits.
  // For now, there is not hardware logic to detect and handle the issue that all the ways in the
  // same set are lock. And it is a programmer's responsibility to make sure that there is at least 
  // one unlock way in a set at any time. 
  // For future backup LRU enhancement project: For pseudo tree LRU algorithm, an efficient backup 
  // LRU algorithm should update the active LRU bits as much as possible, otherwise, it is very possible
  // that the LRU way falls back to the same locked way soon and then forms "LRU trap"
  logic [lg_ways_lp-1:0] lru_way_id;

  logic [ways_p-2:0] modify_mask_lo;
  logic [ways_p-2:0] modify_data_lo;
  logic [ways_p-2:0] modified_lru_bits;

  bsg_lru_pseudo_tree_backup #(
    .ways_p(ways_p)
  ) backup_lru (
    .disabled_ways_i(lock_v_r)
    ,.modify_mask_o(modify_mask_lo)
    ,.modify_data_o(modify_data_lo)
  );

  bsg_mux_bitwise #(
    .width_p(ways_p-1)
  ) lru_bit_mux (
    .data0_i(stat_info_in.lru_bits)
    ,.data1_i(modify_data_lo)
    ,.sel_i(modify_mask_lo)
    ,.data_o(modified_lru_bits)
  );

  bsg_lru_pseudo_tree_encode #(
    .ways_p(ways_p)
  ) lru_encode (
    .lru_i(modified_lru_bits)
    ,.way_id_o(lru_way_id)
  );

  // chosen way demux
  //
  logic [ways_p-1:0] chosen_way_decode;
  bsg_decode #(
    .num_out_p(ways_p)
  ) chosen_way_demux (
    .i(chosen_way_n)
    ,.o(chosen_way_decode)
  );

  // flush way demux
  logic [ways_p-1:0] addr_way_v_r_decode;
  bsg_decode #(
    .num_out_p(ways_p)
  ) addr_way_v_r_demux (
    .i(addr_way_v_r)
    ,.o(addr_way_v_r_decode)
  );
  
  logic [ways_p-1:0] flush_way_decode;
  assign flush_way_decode =  decode_v_r.tagfl_op
    ? addr_way_v_r_decode
    : tag_hit_v_r;

  assign select_snoop_data_r_o = select_snoop_data_r;	

	logic from_evict_data;
	logic from_evict_data_r;

	always_ff @(posedge clk_i) begin
		from_evict_data_r <= from_evict_data;
	end

  always_comb begin

    stat_mem_v_o = 1'b0;
    stat_mem_w_o = 1'b0;
    stat_mem_data_out = '0;
    stat_mem_w_mask_out = '0;

    tag_mem_v_o = 1'b0;
    tag_mem_w_o = 1'b0;
    tag_mem_data_out = '0;
    tag_mem_w_mask_out = '0;

    track_mem_v_o = 1'b0;
    track_mem_w_o = 1'b0;
    track_mem_data_o = '0;
    track_mem_w_mask_o = '0;

    chosen_way_n = chosen_way_r;
    flush_way_n = flush_way_r;

    dma_addr_o = '0;
    dma_cmd_o = e_dma_nop;

    recover_o = '0;
    done_o = '0;

    select_snoop_data_n = select_snoop_data_r;

		miss_state_n = miss_state_r;
		from_evict_data = from_evict_data_r;

    dma_stall_o = 1'b0;

    case (miss_state_r)

      // miss handler waits in this state, until the miss is detected in tv
      // stage.
      // Waits for store buffer and trace buffer to drain then takes over the
      // muxes to the ports to the rams
      START: begin
        // Don't wait for store buffer and trace buffer to drain. Just go.
        //stat_mem_v_o = (miss_v_i & sbuf_empty_i & tbuf_empty_i);
        //track_mem_v_o = word_tracking_p ? (miss_v_i & sbuf_empty_i & tbuf_empty_i) : 1'b0;
        //miss_state_n = (miss_v_i & sbuf_empty_i & tbuf_empty_i)
        //miss_state_n = miss_v ? (goto_flush_op_r ? FLUSH_OP : (goto_lock_op_r ? LOCK_OP 
				//: (st_tag_miss_op_r ? STORE_TAG_MISS : SEND_FILL_ADDR))) : START;

				if(miss_v_i) begin
					if(goto_flush_op_r) begin
						miss_state_n = FLUSH_OP;
					end else if(goto_lock_op_r) begin
						miss_state_n = LOCK_OP;
					end else if(st_tag_miss_op_r) begin
						miss_state_n = STORE_TAG_MISS;
					end else begin
						miss_state_n = SEND_FILL_ADDR;
					end
				end
      end

      // Send out the missing cache block address (to read).
      // Choose a block to replace/fill.
      // If the chosen block is dirty, then take evict route.
      SEND_FILL_ADDR: begin

        // Replacement Policy:
        // If an invalid and unlocked way exists, pick that.
        // If not, pick the LRU way. But if the LRU way designated 
        // by stats_mem_info is locked, it will be overridden by 
        // the bsg_lru_pseudo_tree_backup.
        // On track miss, the chosen way is the tag hit way.
        chosen_way_n = track_miss_r ? tag_hit_way_id_r : (invalid_exist ? invalid_way_id : lru_way_id);

        dma_cmd_o = e_dma_send_fill_addr;
        dma_addr_o = {
          addr_tag_v_r,
          addr_index_v_r,
          {(block_offset_width_lp){1'b0}}
        };

        // if the chosen way is dirty and valid, then evict.
        //miss_state_n = dma_done_i ? ((~track_miss_r & stat_info_in.dirty[chosen_way_n] & valid_v_r[chosen_way_n]) ? SEND_EVICT_ADDR
        //    : GET_FILL_DATA)
        //  : SEND_FILL_ADDR;

        if(dma_done_i) begin
					if(~track_miss_r & stat_info_in.dirty[chosen_way_n] & valid_v_r[chosen_way_n]) begin
						miss_state_n = SEND_EVICT_ADDR;
					end	else begin
						miss_state_n = GET_FILL_DATA;
          end
				end
      end

      // Handling the cases for TAGFL, AINV, AFL, AFLINV.
      FLUSH_OP: begin

        // for TAGFL, pick whichever way set by the addr input.
        // Otherwise, pick the way with the tag hit.
        flush_way_n = decode_v_r.tagfl_op
          ? addr_way_v_r 
          : tag_hit_way_id_r;

        // Clear the dirty bit for the chosen set.
        // LRU bit does not need to be updated.
        stat_mem_v_o = 1'b1;
        stat_mem_w_o = 1'b1;
        stat_mem_data_out.dirty = {ways_p{1'b0}};
        stat_mem_data_out.lru_bits = {(ways_p-1){1'b0}};
        stat_mem_w_mask_out.dirty = flush_way_decode;
        stat_mem_w_mask_out.lru_bits = {(ways_p-1){1'b0}};

        // If it's invalidate op, then clear the valid bit for the chosen way.
        // Otherwise, do not touch the valid bits.
        tag_mem_v_o = 1'b1;
        tag_mem_w_o = 1'b1;

        for (integer i = 0; i < ways_p; i++) begin
          tag_mem_data_out[i].valid = 1'b0;
          tag_mem_data_out[i].lock = 1'b0;
          tag_mem_data_out[i].tag = {tag_width_lp{1'b0}};
          tag_mem_w_mask_out[i].valid = (decode_v_r.ainv_op | decode_v_r.aflinv_op) & flush_way_decode[i];
          tag_mem_w_mask_out[i].lock = (decode_v_r.ainv_op | decode_v_r.aflinv_op) & flush_way_decode[i];
          tag_mem_w_mask_out[i].tag =  {tag_width_lp{1'b0}};
        end

        // If it's not AINV, and the chosen set is dirty and valid, evict the
        // block.
        //miss_state_n = (~decode_v_r.ainv_op & stat_info_in.dirty[flush_way_n] & valid_v_r[flush_way_n])
        //  ? SEND_EVICT_ADDR
        //  : RECOVER;
				if(~decode_v_r.ainv_op & stat_info_in.dirty[flush_way_n] & valid_v_r[flush_way_n]) begin
					miss_state_n = SEND_EVICT_ADDR;
				end else begin
					miss_state_n = RECOVER;
				end
      end

      // handling AUNLOCK, and ALOCK with line not missing.
      LOCK_OP: begin
        tag_mem_v_o = 1'b1;
        tag_mem_w_o = 1'b1;

        for (integer i = 0; i < ways_p; i++) begin
          tag_mem_data_out[i].valid = 1'b0;
          tag_mem_data_out[i].lock = decode_v_r.alock_op;
          tag_mem_data_out[i].tag = {tag_width_lp{1'b0}};
          tag_mem_w_mask_out[i].valid = 1'b0;
          tag_mem_w_mask_out[i].lock = tag_hit_v_r[i];
          tag_mem_w_mask_out[i].tag = {tag_width_lp{1'b0}};
        end
        miss_state_n = RECOVER;
      end

      // Send out the block addr for eviction, before initiating the eviction.
      SEND_EVICT_ADDR: begin
        dma_cmd_o = e_dma_send_evict_addr;
        dma_addr_o = {
          tag_v_r[dma_way_o],
          addr_index_v_r,
          {(block_offset_width_lp){1'b0}}
        };

        //miss_state_n = dma_done_i
        //  ? SEND_EVICT_DATA
        //  : SEND_EVICT_ADDR;
				if(dma_done_i) begin
					miss_state_n = SEND_EVICT_DATA;
				end
      end

      // Set the DMA engine to evict the dirty block.
      // For the flush ops, go straight to RECOVER.
      SEND_EVICT_DATA: begin
        dma_stall_o = 1'b1;
        if(sbuf_empty_i & tbuf_empty_i) begin
            dma_cmd_o = e_dma_send_evict_data;
            dma_addr_o = {
            tag_v_r[dma_way_o],
            addr_index_v_r,
            {(block_offset_width_lp){1'b0}}
          };

          // set stat mem entry on store tag miss.
          stat_mem_v_o = dma_done_i & st_tag_miss_op_r;
          stat_mem_w_o = 1'b1;
          stat_mem_data_out.dirty = {ways_p{1'b1}};
          stat_mem_data_out.lru_bits = chosen_way_lru_data;
          stat_mem_w_mask_out.dirty = chosen_way_decode;
          stat_mem_w_mask_out.lru_bits = chosen_way_lru_mask;

          // set the tag and the valid bit to 1'b1 for the chosen way on store tag miss.
          tag_mem_v_o = dma_done_i & st_tag_miss_op_r;
          tag_mem_w_o = 1'b1;

          for (integer i = 0; i < ways_p; i++) begin
            tag_mem_data_out[i].tag = addr_tag_v_r;
            tag_mem_data_out[i].lock = decode_v_r.alock_op;
            tag_mem_data_out[i].valid = 1'b1;
            tag_mem_w_mask_out[i].tag = {tag_width_lp{chosen_way_decode[i]}};
            tag_mem_w_mask_out[i].lock = chosen_way_decode[i];
            tag_mem_w_mask_out[i].valid = chosen_way_decode[i];
          end

          // set track bits to zero for the chosen way on store tag miss.
          track_mem_v_o = dma_done_i & st_tag_miss_op_r;
          track_mem_w_o = 1'b1;
          for (integer i = 0; i < ways_p; i++) begin
            track_mem_data_o[i] = {block_size_in_words_p{1'b0}};
            track_mem_w_mask_o[i] = {block_size_in_words_p{chosen_way_decode[i]}};
          end

          //miss_state_n = dma_done_i
          //  ? ((decode_v_r.tagfl_op| decode_v_r.aflinv_op| decode_v_r.afl_op | st_tag_miss_op_r) ? RECOVER : GET_FILL_DATA)
          //  : SEND_EVICT_DATA;
				  if(dma_done_i) begin
				    miss_state_n = RECOVER;
				    from_evict_data = 1'b1;
				  //if(decode_v_r.tagfl_op | decode_v_r.aflinv_op | decode_v_r.afl_op | st_tag_miss_op_r) begin
				  //	miss_state_n = RECOVER;
				  //end else begin
				  //	miss_state_n = GET_FILL_DATA;
				  //end
				  end
        end
      end

      // Set the DMA engine to start writing the new block to the data_mem.
      // Do not start until the store buffer is empty.
      GET_FILL_DATA: begin
        dma_cmd_o = e_dma_get_fill_data;
        dma_addr_o = {
          addr_tag_v_r,
          addr_index_v_r,
          {(block_size_in_words_p > 1){addr_block_offset_v_r}}, // used for snoop data in dma.
          {(lg_data_mask_width_lp){1'b0}}
        };
        miss_state_n = WAIT_FOR_FILL_DATA;
      end
      // What is the behavior of the dma_done_i signal?
      // Will need to be high until sbuf and tbuf are empty
      WAIT_FOR_FILL_DATA: begin 
        if(dma_done_i) begin
          dma_stall_o = 1'b1;
          if(sbuf_empty_i & tbuf_empty_i) begin
            // For store tag miss, set the dirty bit for the chosen way.
            // For load tag miss, clear the dirty bit for the chosen way.
            // For track miss, do not touch the dirty bit for the chosen way.
            // Set the lru_bits, so that the chosen way is not the LRU.
            // We are choosing a way to bring in a new block, which is technically
            // the MRU. lru decode unit generates the next state LRU bits, so that
            // the input way is "not" the LRU way.
            stat_mem_v_o = dma_done_i;
            stat_mem_w_o = 1'b1;
            stat_mem_data_out.dirty = {ways_p{decode_v_r.st_op | decode_v_r.atomic_op}};
            stat_mem_data_out.lru_bits = chosen_way_lru_data;
            stat_mem_w_mask_out.dirty = track_miss_r ? {ways_p{1'b0}} : chosen_way_decode;
            stat_mem_w_mask_out.lru_bits = chosen_way_lru_mask;

            // set the tag and the valid bit to 1'b1 for the chosen way.
            tag_mem_v_o = dma_done_i;
            tag_mem_w_o = 1'b1;

            for (integer i = 0; i < ways_p; i++) begin
              tag_mem_data_out[i].tag = addr_tag_v_r;
              tag_mem_data_out[i].lock = decode_v_r.alock_op;
              tag_mem_data_out[i].valid = 1'b1; 
              tag_mem_w_mask_out[i].tag = {tag_width_lp{chosen_way_decode[i]}};
              tag_mem_w_mask_out[i].lock = chosen_way_decode[i];
              tag_mem_w_mask_out[i].valid = chosen_way_decode[i];
            end

            // set track bits to one for the chosen way on store tag miss.
            track_mem_v_o = word_tracking_p ? dma_done_i : 1'b0;
            track_mem_w_o = 1'b1;
            for (integer i = 0; i < ways_p; i++) begin
              track_mem_data_o[i] = {block_size_in_words_p{1'b1}};
              track_mem_w_mask_o[i] = {block_size_in_words_p{chosen_way_decode[i]}};
            end

            select_snoop_data_n = dma_done_i ? 1'b1 : select_snoop_data_r;

            //miss_state_n = dma_done_i
            //  ? RECOVER
            //  : GET_FILL_DATA;
				    if(dma_done_i) begin
				      miss_state_n = RECOVER;
				    end
          end
        end
      end

      // Set the chosen way register. If the line is dirty and valid, evict. 
      // If valid and not dirty, don't evict
      // If not valid, don't evict
      STORE_TAG_MISS: begin
        chosen_way_n = invalid_exist ? invalid_way_id : lru_way_id;

        // if the chosen way is dirty and valid, then evict.
        //miss_state_n = (stat_info_in.dirty[chosen_way_n] & valid_v_r[chosen_way_n])
        //  ? SEND_EVICT_ADDR
        //  : STORE_TAG_MISS_ALLOCATE;
				if(stat_info_in.dirty[chosen_way_n] & valid_v_r[chosen_way_n]) begin
          // Read from the data memory
					miss_state_n = SEND_EVICT_ADDR;
				end else begin
          // Update the tag in the tag memory and write to memory without
          // eviction
					miss_state_n = STORE_TAG_MISS_ALLOCATE;
				end
      end

      STORE_TAG_MISS_ALLOCATE: begin
		    // Write to stat mem
        stat_mem_v_o = 1'b1;
        stat_mem_w_o = 1'b1;
        stat_mem_data_out.dirty = {ways_p{1'b1}};
        stat_mem_data_out.lru_bits = chosen_way_lru_data;
        stat_mem_w_mask_out.dirty = chosen_way_decode;
        stat_mem_w_mask_out.lru_bits = chosen_way_lru_mask;
			
		    // Write to tag mem
        tag_mem_v_o = 1'b1;
        tag_mem_w_o = 1'b1;
        for (integer i = 0; i < ways_p; i++) begin
          tag_mem_data_out[i].tag = addr_tag_v_r;
          tag_mem_data_out[i].lock = decode_v_r.alock_op;
          tag_mem_data_out[i].valid = 1'b1;
          tag_mem_w_mask_out[i].tag = {tag_width_lp{chosen_way_decode[i]}};
          tag_mem_w_mask_out[i].lock = chosen_way_decode[i];
          tag_mem_w_mask_out[i].valid = chosen_way_decode[i];
        end
				
		    // Write to track mem
        track_mem_v_o = 1'b1;
        track_mem_w_o = 1'b1;
        for (integer i = 0; i < ways_p; i++) begin
          track_mem_data_o[i] = {block_size_in_words_p{1'b0}};
          track_mem_w_mask_o[i] = {block_size_in_words_p{chosen_way_decode[i]}};
        end
				
		    // Recover
        miss_state_n = RECOVER;
      end

      // Spend one cycle to recover the tl stage.
      // By recovering, it means re-reading the data_mem and tag_mem for the tl
      // stage.
      RECOVER: begin
        recover_o = 1'b1;
				if(from_evict_data_r) begin
					miss_state_n = GET_FILL_DATA;
					from_evict_data = 1'b0;
				end else begin
        	miss_state_n = DONE;
				end
      end

      // Miss handling is done. Output is valid.
      // Move onto next state, when the output data is taken.
      DONE: begin
        done_o = 1'b1;
        miss_state_n = ack_i ? START : DONE;
        select_snoop_data_n = ack_i ? 1'b0 : select_snoop_data_r;
      end

      // this should never happen, but if it does, go back to START;
      default: begin
        miss_state_n = START;
      end

    endcase
  end

  // synopsys sync_set_reset "reset_i"
  always_ff @ (posedge clk_i) begin
    if (reset_i) begin
      miss_state_r <= START;
      chosen_way_r <= '0;
      flush_way_r <= '0;
      select_snoop_data_r <= 1'b0;
      // added to be a little more X pessimism conservative
      track_data_we_o <= 1'b0;
    end
    else begin
      miss_state_r <= miss_state_n;
      chosen_way_r <= chosen_way_n;
      flush_way_r <= flush_way_n;
      select_snoop_data_r <= select_snoop_data_n;
      track_data_we_o <= track_mem_v_o & ~track_mem_w_o;
    end
  end

endmodule

`BSG_ABSTRACT_MODULE(bsg_cache_miss)
